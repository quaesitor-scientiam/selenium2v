// keys - Set of specific key codes
module keys

pub const null = `\ue000`
pub const cancel = `\ue001`
pub const help = `\ue002`
pub const backspace = `\ue003`
pub const back_space = backspace
pub const tab = `\ue004`
pub const clear = `\ue005`
pub const return_key = `\ue006`
pub const enter = `\ue007`
pub const shift = `\ue008`
pub const left_shift = shift
pub const control = `\ue009`
pub const left_control = control
pub const alt = `\ue00a`
pub const left_alt = alt
pub const pause = `\ue00b`
pub const escape = `\ue00c`
pub const space = `\ue00d`
pub const page_up = `\ue00e`
pub const page_down = `\ue00f`
pub const end = `\ue010`
pub const home = `\ue011`
pub const left = `\ue012`
pub const arrow_left = left
pub const up = `\ue013`
pub const arrow_up = up
pub const right = `\ue014`
pub const arrow_right = right
pub const down = `\ue015`
pub const arrow_down = down
pub const insert = `\ue016`
pub const delete = `\ue017`
pub const semicolon = `\ue018`
pub const equals = `\ue019`

// number pad key codes
pub const numpad0 = `\ue01a`
pub const numpad1 = `\ue01b`
pub const numpad2 = `\ue01c`
pub const numpad3 = `\ue01d`
pub const numpad4 = `\ue01e`
pub const numpad5 = `\ue01f`
pub const numpad6 = `\ue020`
pub const numpad7 = `\ue021`
pub const numpad8 = `\ue022`
pub const numpad9 = `\ue023`
pub const multiply = `\ue024`
pub const add = `\ue025`
pub const separator = `\ue026`
pub const subtract = `\ue027`
pub const decimal = `\ue028`
pub const divide = `\ue029`

// Function key codes
pub const f1 = `\ue031`
pub const f2 = `\ue032`
pub const f3 = `\ue033`
pub const f4 = `\ue034`
pub const f5 = `\ue035`
pub const f6 = `\ue036`
pub const f7 = `\ue037`
pub const f8 = `\ue038`
pub const f9 = `\ue039`
pub const f10 = `\ue03a`
pub const f11 = `\ue03b`
pub const f12 = `\ue03c`

pub const meta = `\ue03d`
pub const command = `\ue03d`
pub const zenkaku_hankaku = `\ue040`
