module common

pub enum WindowTypes {
	tab
	window
}
