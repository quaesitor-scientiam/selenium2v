module remote

pub const remote_commands = {
	'Command.NEW_SESSION':                       ['POST', '/session']
	'Command.QUIT':                              ['DELETE', r'/session/$sessionId']
	'Command.W3C_GET_CURRENT_WINDOW_HANDLE':     ['GET', r'/session/$sessionId/window']
	'Command.W3C_GET_WINDOW_HANDLES':            ['GET', r'/session/$sessionId/handles']
	'Command.GET':                               ['POST', r'/session/$sessionId/url']
	'Command.GO_FORWARD':                        ['POST', r'/session/$sessionId/forward']
	'Command.GO_BACK':                           ['POST', r'/session/$sessionId/back']
	'Command.REFRESH':                           ['POST', r'/session/$sessionId/refresh']
	'Command.W3C_EXECUTE_SCRIPT':                ['POST', r'/session/$sessionId/execute/sync']
	'Command.W3C_EXECUTE_SCRIPT_ASYNC':          ['POST', r'/session/$sessionId/execute/async']
	'Command.GET_CURRENT_URL':                   ['GET', r'/session/$sessionId/url']
	'Command.GET_TITLE':                         ['GET', r'/session/$sessionId/title']
	'Command.GET_PAGE_SOURCE':                   ['GET', r'/session/$sessionId/source']
	'Command.SCREENSHOT':                        ['GET', r'/session/$sessionId/screenshot']
	'Command.ELEMENT_SCREENSHOT':                ['GET', r'/session/$sessionId/element/$id/screenshot']
	'Command.FIND_ELEMENT':                      ['POST', r'/session/$sessionId/element']
	'Command.FIND_ELEMENTS':                     ['POST', r'/session/$sessionId/elements']
	'Command.W3C_GET_ACTIVE_ELEMENT':            ['GET', r'/session/$sessionId/element/active']
	'Command.FIND_CHILD_ELEMENT':                ['POST', r'/session/$sessionId/element/$id/element']
	'Command.FIND_CHILD_ELEMENTS':               ['POST', r'/session/$sessionId/element/$id/elements']
	'Command.CLICK_ELEMENT':                     ['POST', r'/session/$sessionId/element/$id/click']
	'Command.CLEAR_ELEMENT':                     ['POST', r'/session/$sessionId/element/$id/clear']
	'Command.GET_ELEMENT_TEXT':                  ['GET', r'/session/$sessionId/element/$id/text']
	'Command.SEND_KEYS_TO_ELEMENT':              ['POST', r'/session/$sessionId/element/$id/value']
	'Command.GET_ELEMENT_TAG_NAME':              ['GET', r'/session/$sessionId/element/$id/name']
	'Command.IS_ELEMENT_SELECTED':               ['GET', r'/session/$sessionId/element/$id/selected']
	'Command.IS_ELEMENT_ENABLED':                ['GET', r'/session/$sessionId/element/$id/enabled']
	'Command.GET_ELEMENT_RECT':                  ['GET', r'/session/$sessionId/element/$id/rect']
	'Command.GET_ELEMENT_ATTRIBUTE':             ['GET',
		r'/session/$sessionId/element/$id/attribute/$name']
	'Command.GET_ELEMENT_PROPERTY':              ['GET',
		r'/session/$sessionId/element/$id/property/$name']
	'Command.GET_ELEMENT_ARIA_ROLE':             ['GET',
		r'/session/$sessionId/element/$id/computedrole']
	'Command.GET_ELEMENT_ARIA_LABEL':            ['GET',
		r'/session/$sessionId/element/$id/computedlabel']
	'Command.GET_SHADOW_ROOT':                   ['GET', r'/session/$sessionId/element/$id/shadow']
	'Command.FIND_ELEMENT_FROM_SHADOW_ROOT':     ['POST',
		r'/session/$sessionId/shadow/$shadowId/element']
	'Command.FIND_ELEMENTS_FROM_SHADOW_ROOT':    ['POST',
		r'/session/$sessionId/shadow/$shadowId/elements']
	'Command.GET_ALL_COOKIES':                   ['GET', r'/session/$sessionId/cookie']
	'Command.ADD_COOKIE':                        ['POST', r'/session/$sessionId/cookie']
	'Command.GET_COOKIE':                        ['GET', r'/session/$sessionId/cookie/$name']
	'Command.DELETE_ALL_COOKIES':                ['DELETE', r'/session/$sessionId/cookie']
	'Command.DELETE_COOKIE':                     ['DELETE', r'/session/$sessionId/cookie/$name']
	'Command.SWITCH_TO_FRAME':                   ['POST', r'/session/$sessionId/frame']
	'Command.SWITCH_TO_PARENT_FRAME':            ['POST', r'/session/$sessionId/frame/parent']
	'Command.SWITCH_TO_WINDOW':                  ['POST', r'/session/$sessionId/window']
	'Command.NEW_WINDOW':                        ['POST', r'/session/$sessionId/window/new']
	'Command.CLOSE':                             ['DELETE', r'/session/$sessionId/window']
	'Command.GET_ELEMENT_VALUE_OF_CSS_PROPERTY': ['GET',
		r'/session/$sessionId/element/$id/css/$propertyName']
	'Command.EXECUTE_ASYNC_SCRIPT':              ['POST', r'/session/$sessionId/execute_async']
	'Command.SET_TIMEOUTS':                      ['POST', r'/session/$sessionId/timeouts']
	'Command.GET_TIMEOUTS':                      ['GET', r'/session/$sessionId/timeouts']
	'Command.W3C_DISMISS_ALERT':                 ['POST', r'/session/$sessionId/alert/dismiss']
	'Command.W3C_ACCEPT_ALERT':                  ['POST', r'/session/$sessionId/alert/accept']
	'Command.W3C_SET_ALERT_VALUE':               ['POST', r'/session/$sessionId/alert/text']
	'Command.W3C_GET_ALERT_TEXT':                ['GET', r'/session/$sessionId/alert/text']
	'Command.W3C_ACTIONS':                       ['POST', r'/session/$sessionId/actions']
	'Command.W3C_CLEAR_ACTIONS':                 ['DELETE', r'/session/$sessionId/actions']
	'Command.SET_WINDOW_RECT':                   ['POST', r'/session/$sessionId/window/rect']
	'Command.GET_WINDOW_RECT':                   ['GET', r'/session/$sessionId/window/rect']
	'Command.W3C_MAXIMIZE_WINDOW':               ['POST', r'/session/$sessionId/window/maximize']
	'Command.SET_SCREEN_ORIENTATION':            ['POST', r'/session/$sessionId/orientation']
	'Command.GET_SCREEN_ORIENTATION':            ['GET', r'/session/$sessionId/orientation']
	'Command.GET_NETWORK_CONNECTION':            ['GET', r'/session/$sessionId/network_connection']
	'Command.SET_NETWORK_CONNECTION':            ['POST', r'/session/$sessionId/network_connection']
	'Command.GET_LOG':                           ['POST', r'/session/$sessionId/se/log']
	'Command.GET_AVAILABLE_LOG_TYPES':           ['GET', r'/session/$sessionId/se/log/types']
	'Command.CURRENT_CONTEXT_HANDLE':            ['GET', r'/session/$sessionId/context']
	'Command.CONTEXT_HANDLES':                   ['GET', r'/session/$sessionId/contexts']
	'Command.SWITCH_TO_CONTEXT':                 ['POST', r'/session/$sessionId/context']
	'Command.FULLSCREEN_WINDOW':                 ['POST', r'/session/$sessionId/window/fullscreen']
	'Command.MINIMIZE_WINDOW':                   ['POST', r'/session/$sessionId/window/minimize']
	'Command.PRINT_PAGE':                        ['POST', r'/session/$sessionId/print']
	'Command.ADD_VIRTUAL_AUTHENTICATOR':         ['POST',
		r'/session/$sessionId/webauthn/authenticator']
	'Command.REMOVE_VIRTUAL_AUTHENTICATOR':      ['DELETE',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId']
	'Command.ADD_CREDENTIAL':                    ['POST',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId/credential']
	'Command.GET_CREDENTIALS':                   ['GET',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId/credentials']
	'Command.REMOVE_CREDENTIAL':                 ['DELETE',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId/credentials/$credentialId']
	'Command.REMOVE_ALL_CREDENTIALS':            ['DELETE',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId/credentials']
	'Command.SET_USER_VERIFIED':                 ['POST',
		r'/session/$sessionId/webauthn/authenticator/$authenticatorId/uv']
	'Command.UPLOAD_FILE':                       ['POST', r'/session/$sessionId/se/file']
	'Command.GET_DOWNLOADABLE_FILES':            ['GET', r'/session/$sessionId/se/files']
	'Command.DOWNLOAD_FILE':                     ['POST', r'/session/$sessionId/se/files']
	'Command.DELETE_DOWNLOADABLE_FILES':         ['DELETE', r'/session/$sessionId/se/files']
	'Command.GET_FEDCM_TITLE':                   ['GET', r'/session/$sessionId/fedcm/gettitle']
	'Command.GET_FEDCM_DIALOG_TYPE':             ['GET', r'/session/$sessionId/fedcm/getdialogtype']
	'Command.GET_FEDCM_ACCOUNT_LIST':            ['GET', r'/session/$sessionId/fedcm/accountlist']
	'Command.CLICK_FEDCM_DIALOG_BUTTON':         ['POST',
		r'/session/$sessionId/fedcm/clickdialogbutton']
	'Command.CANCEL_FEDCM_DIALOG':               ['POST', r'/session/$sessionId/fedcm/canceldialog']
	'Command.SELECT_FEDCM_ACCOUNT':              ['POST', r'/session/$sessionId/fedcm/selectaccount']
	'Command.SET_FEDCM_DELAY':                   ['POST', r'/session/$sessionId/fedcm/setdelayenabled']
	'Command.RESET_FEDCM_COOLDOWN':              ['POST', r'/session/$sessionId/fedcm/resetcooldown']
}
