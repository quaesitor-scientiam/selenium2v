module chromium

import webdriver.remote { RemoteConnection }

struct ChromiumRemoteConnection {
	RemoteConnection
}
