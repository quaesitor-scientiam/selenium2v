module bidi

import webdriver.remote

pub struct Script {
	// conn 	WebSocketConnection
	log_entry_subscribed bool
}

// fn Script.init(conn WebSocketConnection) Script {
// 	return Script{conn: conn}
// }
