module remote

struct ShadowRoot {
	session int
	id      int
}
