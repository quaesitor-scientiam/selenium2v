module webdriver

import os { File }

pub type SubprocessStdAlias = string | int | f32 | File
