module webdriver

pub const selenium_version = '4.29.0.202501231718'
