module remote

struct Mobile {
}
